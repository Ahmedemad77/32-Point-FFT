
`ifndef FFT_CONFIGRATIONS
`define FFT_CONFIGRATIONS


`define DATA_WIDTH 32
`define ADC_DATA_WIDTH 8 
`define INTEGER 16
`define FRACTION 16
`define CLK_PERIOD 10 


`endif 
