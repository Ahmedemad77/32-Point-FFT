`timescale 1ns / 1ps 

module FFT_32 #(
    parameter
    DATA_WIDTH = 16 , 
    INTEGER = 8, 
	FRACTION = 8,
	ADC_DATA_WIDTH = 8
) (


    input clk,
    input reset,
    input PU_enable,


    input [ADC_DATA_WIDTH-1:0] ADC_in0_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in1_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in2_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in3_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in4_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in5_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in6_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in7_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in8_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in9_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in10_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in11_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in12_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in13_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in14_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in15_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in16_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in17_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in18_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in19_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in20_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in21_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in22_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in23_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in24_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in25_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in26_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in27_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in28_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in29_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in30_real,

    input [ADC_DATA_WIDTH-1:0] ADC_in31_real,


	output [DATA_WIDTH-1:0] FFT_RESULT_0_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_0_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_1_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_1_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_2_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_2_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_3_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_3_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_4_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_4_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_5_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_5_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_6_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_6_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_7_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_7_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_8_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_8_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_9_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_9_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_10_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_10_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_11_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_11_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_12_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_12_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_13_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_13_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_14_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_14_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_15_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_15_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_16_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_16_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_17_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_17_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_18_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_18_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_19_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_19_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_20_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_20_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_21_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_21_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_22_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_22_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_23_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_23_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_24_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_24_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_25_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_25_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_26_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_26_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_27_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_27_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_28_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_28_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_29_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_29_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_30_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_30_imag,

	output [DATA_WIDTH-1:0] FFT_RESULT_31_real,
	output [DATA_WIDTH-1:0] FFT_RESULT_31_imag



);


	wire [DATA_WIDTH-1:0] in0_real;
    wire [DATA_WIDTH-1:0] in1_real;
    wire [DATA_WIDTH-1:0] in2_real;
    wire [DATA_WIDTH-1:0] in3_real;
    wire [DATA_WIDTH-1:0] in4_real;
    wire [DATA_WIDTH-1:0] in5_real;
    wire [DATA_WIDTH-1:0] in6_real;
    wire [DATA_WIDTH-1:0] in7_real;
    wire [DATA_WIDTH-1:0] in8_real;
    wire [DATA_WIDTH-1:0] in9_real;
    wire [DATA_WIDTH-1:0] in10_real;
    wire [DATA_WIDTH-1:0] in11_real;
    wire [DATA_WIDTH-1:0] in12_real;
    wire [DATA_WIDTH-1:0] in13_real;
    wire [DATA_WIDTH-1:0] in14_real;
    wire [DATA_WIDTH-1:0] in15_real;
    wire [DATA_WIDTH-1:0] in16_real;
    wire [DATA_WIDTH-1:0] in17_real;
    wire [DATA_WIDTH-1:0] in18_real;
    wire [DATA_WIDTH-1:0] in19_real;
    wire [DATA_WIDTH-1:0] in20_real;
    wire [DATA_WIDTH-1:0] in21_real;
    wire [DATA_WIDTH-1:0] in22_real;
    wire [DATA_WIDTH-1:0] in23_real;
    wire [DATA_WIDTH-1:0] in24_real;
    wire [DATA_WIDTH-1:0] in25_real;
    wire [DATA_WIDTH-1:0] in26_real;
    wire [DATA_WIDTH-1:0] in27_real;
    wire [DATA_WIDTH-1:0] in28_real;
    wire [DATA_WIDTH-1:0] in29_real;
    wire [DATA_WIDTH-1:0] in30_real;
    wire [DATA_WIDTH-1:0] in31_real;

assign  in0_real = {  { (INTEGER-ADC_DATA_WIDTH) {ADC_in0_real[ADC_DATA_WIDTH-1]}}  ,ADC_in0_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in1_real = {  { (INTEGER-ADC_DATA_WIDTH) {ADC_in1_real[ADC_DATA_WIDTH-1]}}  ,ADC_in1_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in2_real = {  { (INTEGER-ADC_DATA_WIDTH) {ADC_in2_real[ADC_DATA_WIDTH-1]}}  ,ADC_in2_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in3_real = {  { (INTEGER-ADC_DATA_WIDTH) {ADC_in3_real[ADC_DATA_WIDTH-1]}}  ,ADC_in3_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in4_real = {  { (INTEGER-ADC_DATA_WIDTH) {ADC_in4_real[ADC_DATA_WIDTH-1]}}  ,ADC_in4_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in5_real = {  { (INTEGER-ADC_DATA_WIDTH) {ADC_in5_real[ADC_DATA_WIDTH-1]}}  ,ADC_in5_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in6_real = {  { (INTEGER-ADC_DATA_WIDTH) {ADC_in6_real[ADC_DATA_WIDTH-1]}}  ,ADC_in6_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in7_real = {  { (INTEGER-ADC_DATA_WIDTH) {ADC_in7_real[ADC_DATA_WIDTH-1]}}  ,ADC_in7_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in8_real = {  { (INTEGER-ADC_DATA_WIDTH) {ADC_in8_real[ADC_DATA_WIDTH-1]}}  ,ADC_in8_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in9_real = {  { (INTEGER-ADC_DATA_WIDTH) {ADC_in9_real[ADC_DATA_WIDTH-1]}}  ,ADC_in9_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in10_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in10_real[ADC_DATA_WIDTH-1]}}   ,ADC_in10_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in11_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in11_real[ADC_DATA_WIDTH-1]}}   ,ADC_in11_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in12_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in12_real[ADC_DATA_WIDTH-1]}}   ,ADC_in12_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in13_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in13_real[ADC_DATA_WIDTH-1]}}   ,ADC_in13_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in14_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in14_real[ADC_DATA_WIDTH-1]}}   ,ADC_in14_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in15_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in15_real[ADC_DATA_WIDTH-1]}}   ,ADC_in15_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in16_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in16_real[ADC_DATA_WIDTH-1]}}   ,ADC_in16_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in17_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in17_real[ADC_DATA_WIDTH-1]}}   ,ADC_in17_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in18_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in18_real[ADC_DATA_WIDTH-1]}}   ,ADC_in18_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in19_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in19_real[ADC_DATA_WIDTH-1]}}   ,ADC_in19_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in20_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in20_real[ADC_DATA_WIDTH-1]}}   ,ADC_in20_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in21_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in21_real[ADC_DATA_WIDTH-1]}}   ,ADC_in21_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in22_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in22_real[ADC_DATA_WIDTH-1]}}   ,ADC_in22_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in23_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in23_real[ADC_DATA_WIDTH-1]}}   ,ADC_in23_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in24_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in24_real[ADC_DATA_WIDTH-1]}}   ,ADC_in24_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in25_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in25_real[ADC_DATA_WIDTH-1]}}   ,ADC_in25_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in26_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in26_real[ADC_DATA_WIDTH-1]}}   ,ADC_in26_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in27_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in27_real[ADC_DATA_WIDTH-1]}}   ,ADC_in27_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in28_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in28_real[ADC_DATA_WIDTH-1]}}   ,ADC_in28_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in29_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in29_real[ADC_DATA_WIDTH-1]}}   ,ADC_in29_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in30_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in30_real[ADC_DATA_WIDTH-1]}}   ,ADC_in30_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
assign  in31_real = { { (INTEGER-ADC_DATA_WIDTH) {ADC_in31_real[ADC_DATA_WIDTH-1]}}   ,ADC_in31_real , {FRACTION{1'b0}}} ; //Sign Extension And fravtion Filling with zeros 
/////////////////////////////////////////////////////////////////////////////
////////////////////////   Selction Control   ///////////////////////////////
/////////////////////////////////////////////////////////////////////////////

reg [2:0]sel;
always @(posedge clk ) begin
    if (reset) begin
        sel<=3'b000;
    end
    else if (PU_enable) begin
        if (sel==3'b100) begin
           sel <=3'b000; 
        end else begin
            sel <=sel+3'b001;
        end
    end 
end
/////////////////////////////////////////////////////////////////////////////
////////////////////////        Constants       //////////// ////////////////
/////////////////////////////////////////////////////////////////////////////

    wire [DATA_WIDTH-1:0]Constant_W0_real;
    wire [DATA_WIDTH-1:0]Constant_W0_imag;

    wire [DATA_WIDTH-1:0]Constant_W1_real;
    wire [DATA_WIDTH-1:0]Constant_W1_imag;

    wire [DATA_WIDTH-1:0]Constant_W2_real;
    wire [DATA_WIDTH-1:0]Constant_W2_imag;

    wire [DATA_WIDTH-1:0]Constant_W3_real;
    wire [DATA_WIDTH-1:0]Constant_W3_imag;

    wire [DATA_WIDTH-1:0]Constant_W4_real;
    wire [DATA_WIDTH-1:0]Constant_W4_imag;

    wire [DATA_WIDTH-1:0]Constant_W5_real;
    wire [DATA_WIDTH-1:0]Constant_W5_imag;

    wire [DATA_WIDTH-1:0]Constant_W6_real;
    wire [DATA_WIDTH-1:0]Constant_W6_imag;

    wire [DATA_WIDTH-1:0]Constant_W7_real;
    wire [DATA_WIDTH-1:0]Constant_W7_imag;

    wire [DATA_WIDTH-1:0]Constant_W8_real;
    wire [DATA_WIDTH-1:0]Constant_W8_imag;

    wire [DATA_WIDTH-1:0]Constant_W9_real;
    wire [DATA_WIDTH-1:0]Constant_W9_imag;

    wire [DATA_WIDTH-1:0]Constant_W10_real;
    wire [DATA_WIDTH-1:0]Constant_W10_imag;

    wire [DATA_WIDTH-1:0]Constant_W11_real;
    wire [DATA_WIDTH-1:0]Constant_W11_imag;

    wire [DATA_WIDTH-1:0]Constant_W12_real;
    wire [DATA_WIDTH-1:0]Constant_W12_imag;

    wire [DATA_WIDTH-1:0]Constant_W13_real;
    wire [DATA_WIDTH-1:0]Constant_W13_imag;

    wire [DATA_WIDTH-1:0]Constant_W14_real;
    wire [DATA_WIDTH-1:0]Constant_W14_imag;

    wire [DATA_WIDTH-1:0]Constant_W15_real;
    wire [DATA_WIDTH-1:0]Constant_W15_imag;
	/////////////////////////////////////////////////////////////////////////////
	////////////////////////  Constans 32 /16/16 ///////////////////////////////
	/////////////////////////////////////////////////////////////////////////////
//	assign Constant_W0_real  = 16'b0000000100000000;
//    assign Constant_W0_imag  = 16'b0000000000000000;
//    assign Constant_W1_real  = 16'b0000000011111011;
//    assign Constant_W1_imag  = 16'b1111111111001111;
//    assign Constant_W2_real  = 16'b0000000011101100;
//    assign Constant_W2_imag  = 16'b1111111110011111;
//    assign Constant_W3_real  = 16'b0000000011010100;
//    assign Constant_W3_imag  = 16'b1111111101110010;
//    assign Constant_W4_real  = 16'b0000000010110101;
//    assign Constant_W4_imag  = 16'b1111111101001011;
//    assign Constant_W5_real  = 16'b0000000010001110;
//    assign Constant_W5_imag  = 16'b1111111100101100;
//    assign Constant_W6_real  = 16'b0000000001100001;
//    assign Constant_W6_imag  = 16'b1111111100010100;
//    assign Constant_W7_real  = 16'b0000000000110001;
//    assign Constant_W7_imag  = 16'b1111111100000101;
//    assign Constant_W8_real  = 16'b0000000000000000;
//    assign Constant_W8_imag  = 16'b1111111100000000;
//    assign Constant_W9_real  = 16'b1111111111001111;
//    assign Constant_W9_imag  = 16'b1111111100000101;
//    assign Constant_W10_real = 16'b1111111110011111;
//    assign Constant_W10_imag = 16'b1111111100010100;
//    assign Constant_W11_real = 16'b1111111101110010;
//    assign Constant_W11_imag = 16'b1111111100101100;
//    assign Constant_W12_real = 16'b1111111101001011;
//    assign Constant_W12_imag = 16'b1111111101001011;
//    assign Constant_W13_real = 16'b1111111100101100;
//    assign Constant_W13_imag = 16'b1111111101110010;
//    assign Constant_W14_real = 16'b1111111100010100;
//    assign Constant_W14_imag = 16'b1111111110011111;
//    assign Constant_W15_real = 16'b1111111100000101;
//    assign Constant_W15_imag = 16'b1111111111001111;
     assign Constant_W0_real  = 32'b00000000000000010000000000000000;
     assign Constant_W0_imag  = 32'b00000000000000000000000000000000;
     assign Constant_W1_real  = 32'b00000000000000001111101100010100;
     assign Constant_W1_imag  = 32'b11111111111111111100111000001111;
     assign Constant_W2_real  = 32'b00000000000000001110110010000011;
     assign Constant_W2_imag  = 32'b11111111111111111001111000001001;
     assign Constant_W3_real  = 32'b00000000000000001101010011011011;
     assign Constant_W3_imag  = 32'b11111111111111110111000111000111;
     assign Constant_W4_real  = 32'b00000000000000001011010100000100;
     assign Constant_W4_imag  = 32'b11111111111111110100101011111100;
     assign Constant_W5_real  = 32'b00000000000000001000111000111001;
     assign Constant_W5_imag  = 32'b11111111111111110010101100100101;
     assign Constant_W6_real  = 32'b00000000000000000110000111110111;
     assign Constant_W6_imag  = 32'b11111111111111110001001101111101;
     assign Constant_W7_real  = 32'b00000000000000000011000111110001;
     assign Constant_W7_imag  = 32'b11111111111111110000010011101100;
     assign Constant_W8_real  = 32'b00000000000000000000000000000000;
     assign Constant_W8_imag  = 32'b11111111111111110000000000000000;
     assign Constant_W9_real  = 32'b11111111111111111100111000001111;
     assign Constant_W9_imag  = 32'b11111111111111110000010011101100;
     assign Constant_W10_real = 32'b11111111111111111001111000001001;
     assign Constant_W10_imag = 32'b11111111111111110001001101111101;
     assign Constant_W11_real = 32'b11111111111111110111000111000111;
     assign Constant_W11_imag = 32'b11111111111111110010101100100101;
     assign Constant_W12_real = 32'b11111111111111110100101011111100;
     assign Constant_W12_imag = 32'b11111111111111110100101011111100;
     assign Constant_W13_real = 32'b11111111111111110010101100100101;
     assign Constant_W13_imag = 32'b11111111111111110111000111000111;
     assign Constant_W14_real = 32'b11111111111111110001001101111101;
     assign Constant_W14_imag = 32'b11111111111111111001111000001001;
     assign Constant_W15_real = 32'b11111111111111110000010011101100;
     assign Constant_W15_imag = 32'b11111111111111111100111000001111;


/////////////////////////////////////////////////////////////////////////////
////////////////////////        STAGE1       ///////////////////////////////
/////////////////////////////////////////////////////////////////////////////

    wire [DATA_WIDTH-1:0]Stage1_out0_real;
    wire [DATA_WIDTH-1:0]Stage1_out0_imag;
    wire [DATA_WIDTH-1:0]Stage1_out1_real;
    wire [DATA_WIDTH-1:0]Stage1_out1_imag;
    wire [DATA_WIDTH-1:0]Stage1_out2_real;
    wire [DATA_WIDTH-1:0]Stage1_out2_imag;
    wire [DATA_WIDTH-1:0]Stage1_out3_real;
    wire [DATA_WIDTH-1:0]Stage1_out3_imag;
    wire [DATA_WIDTH-1:0]Stage1_out4_real;
    wire [DATA_WIDTH-1:0]Stage1_out4_imag;
    wire [DATA_WIDTH-1:0]Stage1_out5_real;
    wire [DATA_WIDTH-1:0]Stage1_out5_imag;
    wire [DATA_WIDTH-1:0]Stage1_out6_real;
    wire [DATA_WIDTH-1:0]Stage1_out6_imag;
    wire [DATA_WIDTH-1:0]Stage1_out7_real;
    wire [DATA_WIDTH-1:0]Stage1_out7_imag;
    wire [DATA_WIDTH-1:0]Stage1_out8_real;
    wire [DATA_WIDTH-1:0]Stage1_out8_imag;
    wire [DATA_WIDTH-1:0]Stage1_out9_real;
    wire [DATA_WIDTH-1:0]Stage1_out9_imag;
    wire [DATA_WIDTH-1:0]Stage1_out10_real;
    wire [DATA_WIDTH-1:0]Stage1_out10_imag;
    wire [DATA_WIDTH-1:0]Stage1_out11_real;
    wire [DATA_WIDTH-1:0]Stage1_out11_imag;
    wire [DATA_WIDTH-1:0]Stage1_out12_real;
    wire [DATA_WIDTH-1:0]Stage1_out12_imag;
    wire [DATA_WIDTH-1:0]Stage1_out13_real;
    wire [DATA_WIDTH-1:0]Stage1_out13_imag;
    wire [DATA_WIDTH-1:0]Stage1_out14_real;
    wire [DATA_WIDTH-1:0]Stage1_out14_imag;
    wire [DATA_WIDTH-1:0]Stage1_out15_real;
    wire [DATA_WIDTH-1:0]Stage1_out15_imag;
    wire [DATA_WIDTH-1:0]Stage1_out16_real;
    wire [DATA_WIDTH-1:0]Stage1_out16_imag;
    wire [DATA_WIDTH-1:0]Stage1_out17_real;
    wire [DATA_WIDTH-1:0]Stage1_out17_imag;
    wire [DATA_WIDTH-1:0]Stage1_out18_real;
    wire [DATA_WIDTH-1:0]Stage1_out18_imag;
    wire [DATA_WIDTH-1:0]Stage1_out19_real;
    wire [DATA_WIDTH-1:0]Stage1_out19_imag;
    wire [DATA_WIDTH-1:0]Stage1_out20_real;
    wire [DATA_WIDTH-1:0]Stage1_out20_imag;
    wire [DATA_WIDTH-1:0]Stage1_out21_real;
    wire [DATA_WIDTH-1:0]Stage1_out21_imag;
    wire [DATA_WIDTH-1:0]Stage1_out22_real;
    wire [DATA_WIDTH-1:0]Stage1_out22_imag;
    wire [DATA_WIDTH-1:0]Stage1_out23_real;
    wire [DATA_WIDTH-1:0]Stage1_out23_imag;
    wire [DATA_WIDTH-1:0]Stage1_out24_real;
    wire [DATA_WIDTH-1:0]Stage1_out24_imag;
    wire [DATA_WIDTH-1:0]Stage1_out25_real;
    wire [DATA_WIDTH-1:0]Stage1_out25_imag;
    wire [DATA_WIDTH-1:0]Stage1_out26_real;
    wire [DATA_WIDTH-1:0]Stage1_out26_imag;
    wire [DATA_WIDTH-1:0]Stage1_out27_real;
    wire [DATA_WIDTH-1:0]Stage1_out27_imag;
    wire [DATA_WIDTH-1:0]Stage1_out28_real;
    wire [DATA_WIDTH-1:0]Stage1_out28_imag;
    wire [DATA_WIDTH-1:0]Stage1_out29_real;
    wire [DATA_WIDTH-1:0]Stage1_out29_imag;
    wire [DATA_WIDTH-1:0]Stage1_out30_real;
    wire [DATA_WIDTH-1:0]Stage1_out30_imag;
    wire [DATA_WIDTH-1:0]Stage1_out31_real;
    wire [DATA_WIDTH-1:0]Stage1_out31_imag;




FFT_Stage1  #( .DATA_WIDTH(DATA_WIDTH),
.INTEGER(INTEGER),
.FRACTION(FRACTION) ) 

FFT_Stage1Unit (	.clk(clk),
	.reset(reset),
	.PU_enable(PU_enable),
	.sel(sel),
	.in0_real(in0_real),
	.in1_real(in1_real),
	.in2_real(in2_real),
	.in3_real(in3_real),
	.in4_real(in4_real),
	.in5_real(in5_real),
	.in6_real(in6_real),
	.in7_real(in7_real),
	.in8_real(in8_real),
	.in9_real(in9_real),
	.in10_real(in10_real),
	.in11_real(in11_real),
	.in12_real(in12_real),
	.in13_real(in13_real),
	.in14_real(in14_real),
	.in15_real(in15_real),
	.in16_real(in16_real),
	.in17_real(in17_real),
	.in18_real(in18_real),
	.in19_real(in19_real),
	.in20_real(in20_real),
	.in21_real(in21_real),
	.in22_real(in22_real),
	.in23_real(in23_real),
	.in24_real(in24_real),
	.in25_real(in25_real),
	.in26_real(in26_real),
	.in27_real(in27_real),
	.in28_real(in28_real),
	.in29_real(in29_real),
	.in30_real(in30_real),
	.in31_real(in31_real),
	.Constant_W0(Constant_W0_real),
	.Stage1_out0_real(Stage1_out0_real),
	.Stage1_out0_imag(Stage1_out0_imag),
	.Stage1_out1_real(Stage1_out1_real),
	.Stage1_out1_imag(Stage1_out1_imag),
	.Stage1_out2_real(Stage1_out2_real),
	.Stage1_out2_imag(Stage1_out2_imag),
	.Stage1_out3_real(Stage1_out3_real),
	.Stage1_out3_imag(Stage1_out3_imag),
	.Stage1_out4_real(Stage1_out4_real),
	.Stage1_out4_imag(Stage1_out4_imag),
	.Stage1_out5_real(Stage1_out5_real),
	.Stage1_out5_imag(Stage1_out5_imag),
	.Stage1_out6_real(Stage1_out6_real),
	.Stage1_out6_imag(Stage1_out6_imag),
	.Stage1_out7_real(Stage1_out7_real),
	.Stage1_out7_imag(Stage1_out7_imag),
	.Stage1_out8_real(Stage1_out8_real),
	.Stage1_out8_imag(Stage1_out8_imag),
	.Stage1_out9_real(Stage1_out9_real),
	.Stage1_out9_imag(Stage1_out9_imag),
	.Stage1_out10_real(Stage1_out10_real),
	.Stage1_out10_imag(Stage1_out10_imag),
	.Stage1_out11_real(Stage1_out11_real),
	.Stage1_out11_imag(Stage1_out11_imag),
	.Stage1_out12_real(Stage1_out12_real),
	.Stage1_out12_imag(Stage1_out12_imag),
	.Stage1_out13_real(Stage1_out13_real),
	.Stage1_out13_imag(Stage1_out13_imag),
	.Stage1_out14_real(Stage1_out14_real),
	.Stage1_out14_imag(Stage1_out14_imag),
	.Stage1_out15_real(Stage1_out15_real),
	.Stage1_out15_imag(Stage1_out15_imag),
	.Stage1_out16_real(Stage1_out16_real),
	.Stage1_out16_imag(Stage1_out16_imag),
	.Stage1_out17_real(Stage1_out17_real),
	.Stage1_out17_imag(Stage1_out17_imag),
	.Stage1_out18_real(Stage1_out18_real),
	.Stage1_out18_imag(Stage1_out18_imag),
	.Stage1_out19_real(Stage1_out19_real),
	.Stage1_out19_imag(Stage1_out19_imag),
	.Stage1_out20_real(Stage1_out20_real),
	.Stage1_out20_imag(Stage1_out20_imag),
	.Stage1_out21_real(Stage1_out21_real),
	.Stage1_out21_imag(Stage1_out21_imag),
	.Stage1_out22_real(Stage1_out22_real),
	.Stage1_out22_imag(Stage1_out22_imag),
	.Stage1_out23_real(Stage1_out23_real),
	.Stage1_out23_imag(Stage1_out23_imag),
	.Stage1_out24_real(Stage1_out24_real),
	.Stage1_out24_imag(Stage1_out24_imag),
	.Stage1_out25_real(Stage1_out25_real),
	.Stage1_out25_imag(Stage1_out25_imag),
	.Stage1_out26_real(Stage1_out26_real),
	.Stage1_out26_imag(Stage1_out26_imag),
	.Stage1_out27_real(Stage1_out27_real),
	.Stage1_out27_imag(Stage1_out27_imag),
	.Stage1_out28_real(Stage1_out28_real),
	.Stage1_out28_imag(Stage1_out28_imag),
	.Stage1_out29_real(Stage1_out29_real),
	.Stage1_out29_imag(Stage1_out29_imag),
	.Stage1_out30_real(Stage1_out30_real),
	.Stage1_out30_imag(Stage1_out30_imag),
	.Stage1_out31_real(Stage1_out31_real),
	.Stage1_out31_imag(Stage1_out31_imag)
);


/////////////////////////////////////////////////////////////////////////////
////////////////////////        STAGE2       ///////////////////////////////
/////////////////////////////////////////////////////////////////////////////
    wire [DATA_WIDTH-1:0]Stage2_out0_real;
    wire [DATA_WIDTH-1:0]Stage2_out0_imag;
    wire [DATA_WIDTH-1:0]Stage2_out1_real;
    wire [DATA_WIDTH-1:0]Stage2_out1_imag;
    wire [DATA_WIDTH-1:0]Stage2_out2_real;
    wire [DATA_WIDTH-1:0]Stage2_out2_imag;
    wire [DATA_WIDTH-1:0]Stage2_out3_real;
    wire [DATA_WIDTH-1:0]Stage2_out3_imag;
    wire [DATA_WIDTH-1:0]Stage2_out4_real;
    wire [DATA_WIDTH-1:0]Stage2_out4_imag;
    wire [DATA_WIDTH-1:0]Stage2_out5_real;
    wire [DATA_WIDTH-1:0]Stage2_out5_imag;
    wire [DATA_WIDTH-1:0]Stage2_out6_real;
    wire [DATA_WIDTH-1:0]Stage2_out6_imag;
    wire [DATA_WIDTH-1:0]Stage2_out7_real;
    wire [DATA_WIDTH-1:0]Stage2_out7_imag;
    wire [DATA_WIDTH-1:0]Stage2_out8_real;
    wire [DATA_WIDTH-1:0]Stage2_out8_imag;
    wire [DATA_WIDTH-1:0]Stage2_out9_real;
    wire [DATA_WIDTH-1:0]Stage2_out9_imag;
    wire [DATA_WIDTH-1:0]Stage2_out10_real;
    wire [DATA_WIDTH-1:0]Stage2_out10_imag;
    wire [DATA_WIDTH-1:0]Stage2_out11_real;
    wire [DATA_WIDTH-1:0]Stage2_out11_imag;
    wire [DATA_WIDTH-1:0]Stage2_out12_real;
    wire [DATA_WIDTH-1:0]Stage2_out12_imag;
    wire [DATA_WIDTH-1:0]Stage2_out13_real;
    wire [DATA_WIDTH-1:0]Stage2_out13_imag;
    wire [DATA_WIDTH-1:0]Stage2_out14_real;
    wire [DATA_WIDTH-1:0]Stage2_out14_imag;
    wire [DATA_WIDTH-1:0]Stage2_out15_real;
    wire [DATA_WIDTH-1:0]Stage2_out15_imag;
    wire [DATA_WIDTH-1:0]Stage2_out16_real;
    wire [DATA_WIDTH-1:0]Stage2_out16_imag;
    wire [DATA_WIDTH-1:0]Stage2_out17_real;
    wire [DATA_WIDTH-1:0]Stage2_out17_imag;
    wire [DATA_WIDTH-1:0]Stage2_out18_real;
    wire [DATA_WIDTH-1:0]Stage2_out18_imag;
    wire [DATA_WIDTH-1:0]Stage2_out19_real;
    wire [DATA_WIDTH-1:0]Stage2_out19_imag;
    wire [DATA_WIDTH-1:0]Stage2_out20_real;
    wire [DATA_WIDTH-1:0]Stage2_out20_imag;
    wire [DATA_WIDTH-1:0]Stage2_out21_real;
    wire [DATA_WIDTH-1:0]Stage2_out21_imag;
    wire [DATA_WIDTH-1:0]Stage2_out22_real;
    wire [DATA_WIDTH-1:0]Stage2_out22_imag;
    wire [DATA_WIDTH-1:0]Stage2_out23_real;
    wire [DATA_WIDTH-1:0]Stage2_out23_imag;
    wire [DATA_WIDTH-1:0]Stage2_out24_real;
    wire [DATA_WIDTH-1:0]Stage2_out24_imag;
    wire [DATA_WIDTH-1:0]Stage2_out25_real;
    wire [DATA_WIDTH-1:0]Stage2_out25_imag;
    wire [DATA_WIDTH-1:0]Stage2_out26_real;
    wire [DATA_WIDTH-1:0]Stage2_out26_imag;
    wire [DATA_WIDTH-1:0]Stage2_out27_real;
    wire [DATA_WIDTH-1:0]Stage2_out27_imag;
    wire [DATA_WIDTH-1:0]Stage2_out28_real;
    wire [DATA_WIDTH-1:0]Stage2_out28_imag;
    wire [DATA_WIDTH-1:0]Stage2_out29_real;
    wire [DATA_WIDTH-1:0]Stage2_out29_imag;
    wire [DATA_WIDTH-1:0]Stage2_out30_real;
    wire [DATA_WIDTH-1:0]Stage2_out30_imag;
    wire [DATA_WIDTH-1:0]Stage2_out31_real;
    wire [DATA_WIDTH-1:0]Stage2_out31_imag;




FFT_Stage2  #( .DATA_WIDTH(DATA_WIDTH),
.INTEGER(INTEGER),
.FRACTION(FRACTION) ) 

FFT_Stage2Unit (	.clk(clk),
	.reset(reset),
	.PU_enable(PU_enable),
	.sel(sel),
	.Stage1_out0_real(Stage1_out0_real),
	.Stage1_out0_imag(Stage1_out0_imag),
	.Stage1_out1_real(Stage1_out1_real),
	.Stage1_out1_imag(Stage1_out1_imag),
	.Stage1_out2_real(Stage1_out2_real),
	.Stage1_out2_imag(Stage1_out2_imag),
	.Stage1_out3_real(Stage1_out3_real),
	.Stage1_out3_imag(Stage1_out3_imag),
	.Stage1_out4_real(Stage1_out4_real),
	.Stage1_out4_imag(Stage1_out4_imag),
	.Stage1_out5_real(Stage1_out5_real),
	.Stage1_out5_imag(Stage1_out5_imag),
	.Stage1_out6_real(Stage1_out6_real),
	.Stage1_out6_imag(Stage1_out6_imag),
	.Stage1_out7_real(Stage1_out7_real),
	.Stage1_out7_imag(Stage1_out7_imag),
	.Stage1_out8_real(Stage1_out8_real),
	.Stage1_out8_imag(Stage1_out8_imag),
	.Stage1_out9_real(Stage1_out9_real),
	.Stage1_out9_imag(Stage1_out9_imag),
	.Stage1_out10_real(Stage1_out10_real),
	.Stage1_out10_imag(Stage1_out10_imag),
	.Stage1_out11_real(Stage1_out11_real),
	.Stage1_out11_imag(Stage1_out11_imag),
	.Stage1_out12_real(Stage1_out12_real),
	.Stage1_out12_imag(Stage1_out12_imag),
	.Stage1_out13_real(Stage1_out13_real),
	.Stage1_out13_imag(Stage1_out13_imag),
	.Stage1_out14_real(Stage1_out14_real),
	.Stage1_out14_imag(Stage1_out14_imag),
	.Stage1_out15_real(Stage1_out15_real),
	.Stage1_out15_imag(Stage1_out15_imag),
	.Stage1_out16_real(Stage1_out16_real),
	.Stage1_out16_imag(Stage1_out16_imag),
	.Stage1_out17_real(Stage1_out17_real),
	.Stage1_out17_imag(Stage1_out17_imag),
	.Stage1_out18_real(Stage1_out18_real),
	.Stage1_out18_imag(Stage1_out18_imag),
	.Stage1_out19_real(Stage1_out19_real),
	.Stage1_out19_imag(Stage1_out19_imag),
	.Stage1_out20_real(Stage1_out20_real),
	.Stage1_out20_imag(Stage1_out20_imag),
	.Stage1_out21_real(Stage1_out21_real),
	.Stage1_out21_imag(Stage1_out21_imag),
	.Stage1_out22_real(Stage1_out22_real),
	.Stage1_out22_imag(Stage1_out22_imag),
	.Stage1_out23_real(Stage1_out23_real),
	.Stage1_out23_imag(Stage1_out23_imag),
	.Stage1_out24_real(Stage1_out24_real),
	.Stage1_out24_imag(Stage1_out24_imag),
	.Stage1_out25_real(Stage1_out25_real),
	.Stage1_out25_imag(Stage1_out25_imag),
	.Stage1_out26_real(Stage1_out26_real),
	.Stage1_out26_imag(Stage1_out26_imag),
	.Stage1_out27_real(Stage1_out27_real),
	.Stage1_out27_imag(Stage1_out27_imag),
	.Stage1_out28_real(Stage1_out28_real),
	.Stage1_out28_imag(Stage1_out28_imag),
	.Stage1_out29_real(Stage1_out29_real),
	.Stage1_out29_imag(Stage1_out29_imag),
	.Stage1_out30_real(Stage1_out30_real),
	.Stage1_out30_imag(Stage1_out30_imag),
	.Stage1_out31_real(Stage1_out31_real),
	.Stage1_out31_imag(Stage1_out31_imag),
	.Constant_W0_real(Constant_W0_real),
	.Constant_W0_imag(Constant_W0_imag),
	.Constant_W8_real(Constant_W8_real),
	.Constant_W8_imag(Constant_W8_imag),
	.Stage2_out0_real(Stage2_out0_real),
	.Stage2_out0_imag(Stage2_out0_imag),
	.Stage2_out1_real(Stage2_out1_real),
	.Stage2_out1_imag(Stage2_out1_imag),
	.Stage2_out2_real(Stage2_out2_real),
	.Stage2_out2_imag(Stage2_out2_imag),
	.Stage2_out3_real(Stage2_out3_real),
	.Stage2_out3_imag(Stage2_out3_imag),
	.Stage2_out4_real(Stage2_out4_real),
	.Stage2_out4_imag(Stage2_out4_imag),
	.Stage2_out5_real(Stage2_out5_real),
	.Stage2_out5_imag(Stage2_out5_imag),
	.Stage2_out6_real(Stage2_out6_real),
	.Stage2_out6_imag(Stage2_out6_imag),
	.Stage2_out7_real(Stage2_out7_real),
	.Stage2_out7_imag(Stage2_out7_imag),
	.Stage2_out8_real(Stage2_out8_real),
	.Stage2_out8_imag(Stage2_out8_imag),
	.Stage2_out9_real(Stage2_out9_real),
	.Stage2_out9_imag(Stage2_out9_imag),
	.Stage2_out10_real(Stage2_out10_real),
	.Stage2_out10_imag(Stage2_out10_imag),
	.Stage2_out11_real(Stage2_out11_real),
	.Stage2_out11_imag(Stage2_out11_imag),
	.Stage2_out12_real(Stage2_out12_real),
	.Stage2_out12_imag(Stage2_out12_imag),
	.Stage2_out13_real(Stage2_out13_real),
	.Stage2_out13_imag(Stage2_out13_imag),
	.Stage2_out14_real(Stage2_out14_real),
	.Stage2_out14_imag(Stage2_out14_imag),
	.Stage2_out15_real(Stage2_out15_real),
	.Stage2_out15_imag(Stage2_out15_imag),
	.Stage2_out16_real(Stage2_out16_real),
	.Stage2_out16_imag(Stage2_out16_imag),
	.Stage2_out17_real(Stage2_out17_real),
	.Stage2_out17_imag(Stage2_out17_imag),
	.Stage2_out18_real(Stage2_out18_real),
	.Stage2_out18_imag(Stage2_out18_imag),
	.Stage2_out19_real(Stage2_out19_real),
	.Stage2_out19_imag(Stage2_out19_imag),
	.Stage2_out20_real(Stage2_out20_real),
	.Stage2_out20_imag(Stage2_out20_imag),
	.Stage2_out21_real(Stage2_out21_real),
	.Stage2_out21_imag(Stage2_out21_imag),
	.Stage2_out22_real(Stage2_out22_real),
	.Stage2_out22_imag(Stage2_out22_imag),
	.Stage2_out23_real(Stage2_out23_real),
	.Stage2_out23_imag(Stage2_out23_imag),
	.Stage2_out24_real(Stage2_out24_real),
	.Stage2_out24_imag(Stage2_out24_imag),
	.Stage2_out25_real(Stage2_out25_real),
	.Stage2_out25_imag(Stage2_out25_imag),
	.Stage2_out26_real(Stage2_out26_real),
	.Stage2_out26_imag(Stage2_out26_imag),
	.Stage2_out27_real(Stage2_out27_real),
	.Stage2_out27_imag(Stage2_out27_imag),
	.Stage2_out28_real(Stage2_out28_real),
	.Stage2_out28_imag(Stage2_out28_imag),
	.Stage2_out29_real(Stage2_out29_real),
	.Stage2_out29_imag(Stage2_out29_imag),
	.Stage2_out30_real(Stage2_out30_real),
	.Stage2_out30_imag(Stage2_out30_imag),
	.Stage2_out31_real(Stage2_out31_real),
	.Stage2_out31_imag(Stage2_out31_imag)
);


/////////////////////////////////////////////////////////////////////////////
////////////////////////        STAGE3       ///////////////////////////////
/////////////////////////////////////////////////////////////////////////////
    wire [DATA_WIDTH-1:0]Stage3_out0_real;
    wire [DATA_WIDTH-1:0]Stage3_out0_imag;
    wire [DATA_WIDTH-1:0]Stage3_out1_real;
    wire [DATA_WIDTH-1:0]Stage3_out1_imag;
    wire [DATA_WIDTH-1:0]Stage3_out2_real;
    wire [DATA_WIDTH-1:0]Stage3_out2_imag;
    wire [DATA_WIDTH-1:0]Stage3_out3_real;
    wire [DATA_WIDTH-1:0]Stage3_out3_imag;
    wire [DATA_WIDTH-1:0]Stage3_out4_real;
    wire [DATA_WIDTH-1:0]Stage3_out4_imag;
    wire [DATA_WIDTH-1:0]Stage3_out5_real;
    wire [DATA_WIDTH-1:0]Stage3_out5_imag;
    wire [DATA_WIDTH-1:0]Stage3_out6_real;
    wire [DATA_WIDTH-1:0]Stage3_out6_imag;
    wire [DATA_WIDTH-1:0]Stage3_out7_real;
    wire [DATA_WIDTH-1:0]Stage3_out7_imag;
    wire [DATA_WIDTH-1:0]Stage3_out8_real;
    wire [DATA_WIDTH-1:0]Stage3_out8_imag;
    wire [DATA_WIDTH-1:0]Stage3_out9_real;
    wire [DATA_WIDTH-1:0]Stage3_out9_imag;
    wire [DATA_WIDTH-1:0]Stage3_out10_real;
    wire [DATA_WIDTH-1:0]Stage3_out10_imag;
    wire [DATA_WIDTH-1:0]Stage3_out11_real;
    wire [DATA_WIDTH-1:0]Stage3_out11_imag;
    wire [DATA_WIDTH-1:0]Stage3_out12_real;
    wire [DATA_WIDTH-1:0]Stage3_out12_imag;
    wire [DATA_WIDTH-1:0]Stage3_out13_real;
    wire [DATA_WIDTH-1:0]Stage3_out13_imag;
    wire [DATA_WIDTH-1:0]Stage3_out14_real;
    wire [DATA_WIDTH-1:0]Stage3_out14_imag;
    wire [DATA_WIDTH-1:0]Stage3_out15_real;
    wire [DATA_WIDTH-1:0]Stage3_out15_imag;
    wire [DATA_WIDTH-1:0]Stage3_out16_real;
    wire [DATA_WIDTH-1:0]Stage3_out16_imag;
    wire [DATA_WIDTH-1:0]Stage3_out17_real;
    wire [DATA_WIDTH-1:0]Stage3_out17_imag;
    wire [DATA_WIDTH-1:0]Stage3_out18_real;
    wire [DATA_WIDTH-1:0]Stage3_out18_imag;
    wire [DATA_WIDTH-1:0]Stage3_out19_real;
    wire [DATA_WIDTH-1:0]Stage3_out19_imag;
    wire [DATA_WIDTH-1:0]Stage3_out20_real;
    wire [DATA_WIDTH-1:0]Stage3_out20_imag;
    wire [DATA_WIDTH-1:0]Stage3_out21_real;
    wire [DATA_WIDTH-1:0]Stage3_out21_imag;
    wire [DATA_WIDTH-1:0]Stage3_out22_real;
    wire [DATA_WIDTH-1:0]Stage3_out22_imag;
    wire [DATA_WIDTH-1:0]Stage3_out23_real;
    wire [DATA_WIDTH-1:0]Stage3_out23_imag;
    wire [DATA_WIDTH-1:0]Stage3_out24_real;
    wire [DATA_WIDTH-1:0]Stage3_out24_imag;
    wire [DATA_WIDTH-1:0]Stage3_out25_real;
    wire [DATA_WIDTH-1:0]Stage3_out25_imag;
    wire [DATA_WIDTH-1:0]Stage3_out26_real;
    wire [DATA_WIDTH-1:0]Stage3_out26_imag;
    wire [DATA_WIDTH-1:0]Stage3_out27_real;
    wire [DATA_WIDTH-1:0]Stage3_out27_imag;
    wire [DATA_WIDTH-1:0]Stage3_out28_real;
    wire [DATA_WIDTH-1:0]Stage3_out28_imag;
    wire [DATA_WIDTH-1:0]Stage3_out29_real;
    wire [DATA_WIDTH-1:0]Stage3_out29_imag;
    wire [DATA_WIDTH-1:0]Stage3_out30_real;
    wire [DATA_WIDTH-1:0]Stage3_out30_imag;
    wire [DATA_WIDTH-1:0]Stage3_out31_real;
    wire [DATA_WIDTH-1:0]Stage3_out31_imag;




FFT_Stage3  #( .DATA_WIDTH(DATA_WIDTH),
.INTEGER(INTEGER),
.FRACTION(FRACTION) ) 

FFT_Stage3Unit (	.clk(clk),
	.reset(reset),
	.PU_enable(PU_enable),
	.sel(sel),
	.Stage2_out0_real(Stage2_out0_real),
	.Stage2_out0_imag(Stage2_out0_imag),
	.Stage2_out1_real(Stage2_out1_real),
	.Stage2_out1_imag(Stage2_out1_imag),
	.Stage2_out2_real(Stage2_out2_real),
	.Stage2_out2_imag(Stage2_out2_imag),
	.Stage2_out3_real(Stage2_out3_real),
	.Stage2_out3_imag(Stage2_out3_imag),
	.Stage2_out4_real(Stage2_out4_real),
	.Stage2_out4_imag(Stage2_out4_imag),
	.Stage2_out5_real(Stage2_out5_real),
	.Stage2_out5_imag(Stage2_out5_imag),
	.Stage2_out6_real(Stage2_out6_real),
	.Stage2_out6_imag(Stage2_out6_imag),
	.Stage2_out7_real(Stage2_out7_real),
	.Stage2_out7_imag(Stage2_out7_imag),
	.Stage2_out8_real(Stage2_out8_real),
	.Stage2_out8_imag(Stage2_out8_imag),
	.Stage2_out9_real(Stage2_out9_real),
	.Stage2_out9_imag(Stage2_out9_imag),
	.Stage2_out10_real(Stage2_out10_real),
	.Stage2_out10_imag(Stage2_out10_imag),
	.Stage2_out11_real(Stage2_out11_real),
	.Stage2_out11_imag(Stage2_out11_imag),
	.Stage2_out12_real(Stage2_out12_real),
	.Stage2_out12_imag(Stage2_out12_imag),
	.Stage2_out13_real(Stage2_out13_real),
	.Stage2_out13_imag(Stage2_out13_imag),
	.Stage2_out14_real(Stage2_out14_real),
	.Stage2_out14_imag(Stage2_out14_imag),
	.Stage2_out15_real(Stage2_out15_real),
	.Stage2_out15_imag(Stage2_out15_imag),
	.Stage2_out16_real(Stage2_out16_real),
	.Stage2_out16_imag(Stage2_out16_imag),
	.Stage2_out17_real(Stage2_out17_real),
	.Stage2_out17_imag(Stage2_out17_imag),
	.Stage2_out18_real(Stage2_out18_real),
	.Stage2_out18_imag(Stage2_out18_imag),
	.Stage2_out19_real(Stage2_out19_real),
	.Stage2_out19_imag(Stage2_out19_imag),
	.Stage2_out20_real(Stage2_out20_real),
	.Stage2_out20_imag(Stage2_out20_imag),
	.Stage2_out21_real(Stage2_out21_real),
	.Stage2_out21_imag(Stage2_out21_imag),
	.Stage2_out22_real(Stage2_out22_real),
	.Stage2_out22_imag(Stage2_out22_imag),
	.Stage2_out23_real(Stage2_out23_real),
	.Stage2_out23_imag(Stage2_out23_imag),
	.Stage2_out24_real(Stage2_out24_real),
	.Stage2_out24_imag(Stage2_out24_imag),
	.Stage2_out25_real(Stage2_out25_real),
	.Stage2_out25_imag(Stage2_out25_imag),
	.Stage2_out26_real(Stage2_out26_real),
	.Stage2_out26_imag(Stage2_out26_imag),
	.Stage2_out27_real(Stage2_out27_real),
	.Stage2_out27_imag(Stage2_out27_imag),
	.Stage2_out28_real(Stage2_out28_real),
	.Stage2_out28_imag(Stage2_out28_imag),
	.Stage2_out29_real(Stage2_out29_real),
	.Stage2_out29_imag(Stage2_out29_imag),
	.Stage2_out30_real(Stage2_out30_real),
	.Stage2_out30_imag(Stage2_out30_imag),
	.Stage2_out31_real(Stage2_out31_real),
	.Stage2_out31_imag(Stage2_out31_imag),
	.Stage3_out0_real(Stage3_out0_real),
	.Stage3_out0_imag(Stage3_out0_imag),
	.Stage3_out1_real(Stage3_out1_real),
	.Stage3_out1_imag(Stage3_out1_imag),
	.Stage3_out2_real(Stage3_out2_real),
	.Stage3_out2_imag(Stage3_out2_imag),
	.Stage3_out3_real(Stage3_out3_real),
	.Stage3_out3_imag(Stage3_out3_imag),
	.Stage3_out4_real(Stage3_out4_real),
	.Stage3_out4_imag(Stage3_out4_imag),
	.Stage3_out5_real(Stage3_out5_real),
	.Stage3_out5_imag(Stage3_out5_imag),
	.Stage3_out6_real(Stage3_out6_real),
	.Stage3_out6_imag(Stage3_out6_imag),
	.Stage3_out7_real(Stage3_out7_real),
	.Stage3_out7_imag(Stage3_out7_imag),
	.Stage3_out8_real(Stage3_out8_real),
	.Stage3_out8_imag(Stage3_out8_imag),
	.Stage3_out9_real(Stage3_out9_real),
	.Stage3_out9_imag(Stage3_out9_imag),
	.Stage3_out10_real(Stage3_out10_real),
	.Stage3_out10_imag(Stage3_out10_imag),
	.Stage3_out11_real(Stage3_out11_real),
	.Stage3_out11_imag(Stage3_out11_imag),
	.Stage3_out12_real(Stage3_out12_real),
	.Stage3_out12_imag(Stage3_out12_imag),
	.Stage3_out13_real(Stage3_out13_real),
	.Stage3_out13_imag(Stage3_out13_imag),
	.Stage3_out14_real(Stage3_out14_real),
	.Stage3_out14_imag(Stage3_out14_imag),
	.Stage3_out15_real(Stage3_out15_real),
	.Stage3_out15_imag(Stage3_out15_imag),
	.Stage3_out16_real(Stage3_out16_real),
	.Stage3_out16_imag(Stage3_out16_imag),
	.Stage3_out17_real(Stage3_out17_real),
	.Stage3_out17_imag(Stage3_out17_imag),
	.Stage3_out18_real(Stage3_out18_real),
	.Stage3_out18_imag(Stage3_out18_imag),
	.Stage3_out19_real(Stage3_out19_real),
	.Stage3_out19_imag(Stage3_out19_imag),
	.Stage3_out20_real(Stage3_out20_real),
	.Stage3_out20_imag(Stage3_out20_imag),
	.Stage3_out21_real(Stage3_out21_real),
	.Stage3_out21_imag(Stage3_out21_imag),
	.Stage3_out22_real(Stage3_out22_real),
	.Stage3_out22_imag(Stage3_out22_imag),
	.Stage3_out23_real(Stage3_out23_real),
	.Stage3_out23_imag(Stage3_out23_imag),
	.Stage3_out24_real(Stage3_out24_real),
	.Stage3_out24_imag(Stage3_out24_imag),
	.Stage3_out25_real(Stage3_out25_real),
	.Stage3_out25_imag(Stage3_out25_imag),
	.Stage3_out26_real(Stage3_out26_real),
	.Stage3_out26_imag(Stage3_out26_imag),
	.Stage3_out27_real(Stage3_out27_real),
	.Stage3_out27_imag(Stage3_out27_imag),
	.Stage3_out28_real(Stage3_out28_real),
	.Stage3_out28_imag(Stage3_out28_imag),
	.Stage3_out29_real(Stage3_out29_real),
	.Stage3_out29_imag(Stage3_out29_imag),
	.Stage3_out30_real(Stage3_out30_real),
	.Stage3_out30_imag(Stage3_out30_imag),
	.Stage3_out31_real(Stage3_out31_real),
	.Stage3_out31_imag(Stage3_out31_imag),
	.Constant_W0_real(Constant_W0_real),
	.Constant_W0_imag(Constant_W0_imag),
	.Constant_W4_real(Constant_W4_real),
	.Constant_W4_imag(Constant_W4_imag),
	.Constant_W8_real(Constant_W8_real),
	.Constant_W8_imag(Constant_W8_imag),
	.Constant_W12_real(Constant_W12_real),
	.Constant_W12_imag(Constant_W12_imag)
);


/////////////////////////////////////////////////////////////////////////////
////////////////////////        STAGE4       ///////////////////////////////
/////////////////////////////////////////////////////////////////////////////
    wire [DATA_WIDTH-1:0]Stage4_out0_real;
    wire [DATA_WIDTH-1:0]Stage4_out0_imag;
    wire [DATA_WIDTH-1:0]Stage4_out1_real;
    wire [DATA_WIDTH-1:0]Stage4_out1_imag;
    wire [DATA_WIDTH-1:0]Stage4_out2_real;
    wire [DATA_WIDTH-1:0]Stage4_out2_imag;
    wire [DATA_WIDTH-1:0]Stage4_out3_real;
    wire [DATA_WIDTH-1:0]Stage4_out3_imag;
    wire [DATA_WIDTH-1:0]Stage4_out4_real;
    wire [DATA_WIDTH-1:0]Stage4_out4_imag;
    wire [DATA_WIDTH-1:0]Stage4_out5_real;
    wire [DATA_WIDTH-1:0]Stage4_out5_imag;
    wire [DATA_WIDTH-1:0]Stage4_out6_real;
    wire [DATA_WIDTH-1:0]Stage4_out6_imag;
    wire [DATA_WIDTH-1:0]Stage4_out7_real;
    wire [DATA_WIDTH-1:0]Stage4_out7_imag;
    wire [DATA_WIDTH-1:0]Stage4_out8_real;
    wire [DATA_WIDTH-1:0]Stage4_out8_imag;
    wire [DATA_WIDTH-1:0]Stage4_out9_real;
    wire [DATA_WIDTH-1:0]Stage4_out9_imag;
    wire [DATA_WIDTH-1:0]Stage4_out10_real;
    wire [DATA_WIDTH-1:0]Stage4_out10_imag;
    wire [DATA_WIDTH-1:0]Stage4_out11_real;
    wire [DATA_WIDTH-1:0]Stage4_out11_imag;
    wire [DATA_WIDTH-1:0]Stage4_out12_real;
    wire [DATA_WIDTH-1:0]Stage4_out12_imag;
    wire [DATA_WIDTH-1:0]Stage4_out13_real;
    wire [DATA_WIDTH-1:0]Stage4_out13_imag;
    wire [DATA_WIDTH-1:0]Stage4_out14_real;
    wire [DATA_WIDTH-1:0]Stage4_out14_imag;
    wire [DATA_WIDTH-1:0]Stage4_out15_real;
    wire [DATA_WIDTH-1:0]Stage4_out15_imag;
    wire [DATA_WIDTH-1:0]Stage4_out16_real;
    wire [DATA_WIDTH-1:0]Stage4_out16_imag;
    wire [DATA_WIDTH-1:0]Stage4_out17_real;
    wire [DATA_WIDTH-1:0]Stage4_out17_imag;
    wire [DATA_WIDTH-1:0]Stage4_out18_real;
    wire [DATA_WIDTH-1:0]Stage4_out18_imag;
    wire [DATA_WIDTH-1:0]Stage4_out19_real;
    wire [DATA_WIDTH-1:0]Stage4_out19_imag;
    wire [DATA_WIDTH-1:0]Stage4_out20_real;
    wire [DATA_WIDTH-1:0]Stage4_out20_imag;
    wire [DATA_WIDTH-1:0]Stage4_out21_real;
    wire [DATA_WIDTH-1:0]Stage4_out21_imag;
    wire [DATA_WIDTH-1:0]Stage4_out22_real;
    wire [DATA_WIDTH-1:0]Stage4_out22_imag;
    wire [DATA_WIDTH-1:0]Stage4_out23_real;
    wire [DATA_WIDTH-1:0]Stage4_out23_imag;
    wire [DATA_WIDTH-1:0]Stage4_out24_real;
    wire [DATA_WIDTH-1:0]Stage4_out24_imag;
    wire [DATA_WIDTH-1:0]Stage4_out25_real;
    wire [DATA_WIDTH-1:0]Stage4_out25_imag;
    wire [DATA_WIDTH-1:0]Stage4_out26_real;
    wire [DATA_WIDTH-1:0]Stage4_out26_imag;
    wire [DATA_WIDTH-1:0]Stage4_out27_real;
    wire [DATA_WIDTH-1:0]Stage4_out27_imag;
    wire [DATA_WIDTH-1:0]Stage4_out28_real;
    wire [DATA_WIDTH-1:0]Stage4_out28_imag;
    wire [DATA_WIDTH-1:0]Stage4_out29_real;
    wire [DATA_WIDTH-1:0]Stage4_out29_imag;
    wire [DATA_WIDTH-1:0]Stage4_out30_real;
    wire [DATA_WIDTH-1:0]Stage4_out30_imag;
    wire [DATA_WIDTH-1:0]Stage4_out31_real;
    wire [DATA_WIDTH-1:0]Stage4_out31_imag;

FFT_Stage4  #( .DATA_WIDTH(DATA_WIDTH),
.INTEGER(INTEGER),
.FRACTION(FRACTION) ) 

FFT_Stage4Unit (	.clk(clk),
	.reset(reset),
	.PU_enable(PU_enable),
	.sel(sel),
	.Stage3_out0_real(Stage3_out0_real),
	.Stage3_out0_imag(Stage3_out0_imag),
	.Stage3_out1_real(Stage3_out1_real),
	.Stage3_out1_imag(Stage3_out1_imag),
	.Stage3_out2_real(Stage3_out2_real),
	.Stage3_out2_imag(Stage3_out2_imag),
	.Stage3_out3_real(Stage3_out3_real),
	.Stage3_out3_imag(Stage3_out3_imag),
	.Stage3_out4_real(Stage3_out4_real),
	.Stage3_out4_imag(Stage3_out4_imag),
	.Stage3_out5_real(Stage3_out5_real),
	.Stage3_out5_imag(Stage3_out5_imag),
	.Stage3_out6_real(Stage3_out6_real),
	.Stage3_out6_imag(Stage3_out6_imag),
	.Stage3_out7_real(Stage3_out7_real),
	.Stage3_out7_imag(Stage3_out7_imag),
	.Stage3_out8_real(Stage3_out8_real),
	.Stage3_out8_imag(Stage3_out8_imag),
	.Stage3_out9_real(Stage3_out9_real),
	.Stage3_out9_imag(Stage3_out9_imag),
	.Stage3_out10_real(Stage3_out10_real),
	.Stage3_out10_imag(Stage3_out10_imag),
	.Stage3_out11_real(Stage3_out11_real),
	.Stage3_out11_imag(Stage3_out11_imag),
	.Stage3_out12_real(Stage3_out12_real),
	.Stage3_out12_imag(Stage3_out12_imag),
	.Stage3_out13_real(Stage3_out13_real),
	.Stage3_out13_imag(Stage3_out13_imag),
	.Stage3_out14_real(Stage3_out14_real),
	.Stage3_out14_imag(Stage3_out14_imag),
	.Stage3_out15_real(Stage3_out15_real),
	.Stage3_out15_imag(Stage3_out15_imag),
	.Stage3_out16_real(Stage3_out16_real),
	.Stage3_out16_imag(Stage3_out16_imag),
	.Stage3_out17_real(Stage3_out17_real),
	.Stage3_out17_imag(Stage3_out17_imag),
	.Stage3_out18_real(Stage3_out18_real),
	.Stage3_out18_imag(Stage3_out18_imag),
	.Stage3_out19_real(Stage3_out19_real),
	.Stage3_out19_imag(Stage3_out19_imag),
	.Stage3_out20_real(Stage3_out20_real),
	.Stage3_out20_imag(Stage3_out20_imag),
	.Stage3_out21_real(Stage3_out21_real),
	.Stage3_out21_imag(Stage3_out21_imag),
	.Stage3_out22_real(Stage3_out22_real),
	.Stage3_out22_imag(Stage3_out22_imag),
	.Stage3_out23_real(Stage3_out23_real),
	.Stage3_out23_imag(Stage3_out23_imag),
	.Stage3_out24_real(Stage3_out24_real),
	.Stage3_out24_imag(Stage3_out24_imag),
	.Stage3_out25_real(Stage3_out25_real),
	.Stage3_out25_imag(Stage3_out25_imag),
	.Stage3_out26_real(Stage3_out26_real),
	.Stage3_out26_imag(Stage3_out26_imag),
	.Stage3_out27_real(Stage3_out27_real),
	.Stage3_out27_imag(Stage3_out27_imag),
	.Stage3_out28_real(Stage3_out28_real),
	.Stage3_out28_imag(Stage3_out28_imag),
	.Stage3_out29_real(Stage3_out29_real),
	.Stage3_out29_imag(Stage3_out29_imag),
	.Stage3_out30_real(Stage3_out30_real),
	.Stage3_out30_imag(Stage3_out30_imag),
	.Stage3_out31_real(Stage3_out31_real),
	.Stage3_out31_imag(Stage3_out31_imag),
	.Stage4_out0_real(Stage4_out0_real),
	.Stage4_out0_imag(Stage4_out0_imag),
	.Stage4_out1_real(Stage4_out1_real),
	.Stage4_out1_imag(Stage4_out1_imag),
	.Stage4_out2_real(Stage4_out2_real),
	.Stage4_out2_imag(Stage4_out2_imag),
	.Stage4_out3_real(Stage4_out3_real),
	.Stage4_out3_imag(Stage4_out3_imag),
	.Stage4_out4_real(Stage4_out4_real),
	.Stage4_out4_imag(Stage4_out4_imag),
	.Stage4_out5_real(Stage4_out5_real),
	.Stage4_out5_imag(Stage4_out5_imag),
	.Stage4_out6_real(Stage4_out6_real),
	.Stage4_out6_imag(Stage4_out6_imag),
	.Stage4_out7_real(Stage4_out7_real),
	.Stage4_out7_imag(Stage4_out7_imag),
	.Stage4_out8_real(Stage4_out8_real),
	.Stage4_out8_imag(Stage4_out8_imag),
	.Stage4_out9_real(Stage4_out9_real),
	.Stage4_out9_imag(Stage4_out9_imag),
	.Stage4_out10_real(Stage4_out10_real),
	.Stage4_out10_imag(Stage4_out10_imag),
	.Stage4_out11_real(Stage4_out11_real),
	.Stage4_out11_imag(Stage4_out11_imag),
	.Stage4_out12_real(Stage4_out12_real),
	.Stage4_out12_imag(Stage4_out12_imag),
	.Stage4_out13_real(Stage4_out13_real),
	.Stage4_out13_imag(Stage4_out13_imag),
	.Stage4_out14_real(Stage4_out14_real),
	.Stage4_out14_imag(Stage4_out14_imag),
	.Stage4_out15_real(Stage4_out15_real),
	.Stage4_out15_imag(Stage4_out15_imag),
	.Stage4_out16_real(Stage4_out16_real),
	.Stage4_out16_imag(Stage4_out16_imag),
	.Stage4_out17_real(Stage4_out17_real),
	.Stage4_out17_imag(Stage4_out17_imag),
	.Stage4_out18_real(Stage4_out18_real),
	.Stage4_out18_imag(Stage4_out18_imag),
	.Stage4_out19_real(Stage4_out19_real),
	.Stage4_out19_imag(Stage4_out19_imag),
	.Stage4_out20_real(Stage4_out20_real),
	.Stage4_out20_imag(Stage4_out20_imag),
	.Stage4_out21_real(Stage4_out21_real),
	.Stage4_out21_imag(Stage4_out21_imag),
	.Stage4_out22_real(Stage4_out22_real),
	.Stage4_out22_imag(Stage4_out22_imag),
	.Stage4_out23_real(Stage4_out23_real),
	.Stage4_out23_imag(Stage4_out23_imag),
	.Stage4_out24_real(Stage4_out24_real),
	.Stage4_out24_imag(Stage4_out24_imag),
	.Stage4_out25_real(Stage4_out25_real),
	.Stage4_out25_imag(Stage4_out25_imag),
	.Stage4_out26_real(Stage4_out26_real),
	.Stage4_out26_imag(Stage4_out26_imag),
	.Stage4_out27_real(Stage4_out27_real),
	.Stage4_out27_imag(Stage4_out27_imag),
	.Stage4_out28_real(Stage4_out28_real),
	.Stage4_out28_imag(Stage4_out28_imag),
	.Stage4_out29_real(Stage4_out29_real),
	.Stage4_out29_imag(Stage4_out29_imag),
	.Stage4_out30_real(Stage4_out30_real),
	.Stage4_out30_imag(Stage4_out30_imag),
	.Stage4_out31_real(Stage4_out31_real),
	.Stage4_out31_imag(Stage4_out31_imag),
	.Constant_W0_real(Constant_W0_real),
	.Constant_W0_imag(Constant_W0_imag),
	.Constant_W2_real(Constant_W2_real),
	.Constant_W2_imag(Constant_W2_imag),
	.Constant_W4_real(Constant_W4_real),
	.Constant_W4_imag(Constant_W4_imag),
	.Constant_W6_real(Constant_W6_real),
	.Constant_W6_imag(Constant_W6_imag),
	.Constant_W8_real(Constant_W8_real),
	.Constant_W8_imag(Constant_W8_imag),
	.Constant_W10_real(Constant_W10_real),
	.Constant_W10_imag(Constant_W10_imag),
	.Constant_W12_real(Constant_W12_real),
	.Constant_W12_imag(Constant_W12_imag),
	.Constant_W14_real(Constant_W14_real),
	.Constant_W14_imag(Constant_W14_imag)
);



/////////////////////////////////////////////////////////////////////////////
////////////////////////        STAGE5        ///////////////////////////////
/////////////////////////////////////////////////////////////////////////////


FFT_Stage5  #( .DATA_WIDTH(DATA_WIDTH),
.INTEGER(INTEGER),
.FRACTION(FRACTION) ) 

FFT_Stage5Unit (	.clk(clk),
	.reset(reset),
	.PU_enable(PU_enable),
	.sel(sel),
	.Stage4_out0_real(Stage4_out0_real),
	.Stage4_out0_imag(Stage4_out0_imag),
	.Stage4_out1_real(Stage4_out1_real),
	.Stage4_out1_imag(Stage4_out1_imag),
	.Stage4_out2_real(Stage4_out2_real),
	.Stage4_out2_imag(Stage4_out2_imag),
	.Stage4_out3_real(Stage4_out3_real),
	.Stage4_out3_imag(Stage4_out3_imag),
	.Stage4_out4_real(Stage4_out4_real),
	.Stage4_out4_imag(Stage4_out4_imag),
	.Stage4_out5_real(Stage4_out5_real),
	.Stage4_out5_imag(Stage4_out5_imag),
	.Stage4_out6_real(Stage4_out6_real),
	.Stage4_out6_imag(Stage4_out6_imag),
	.Stage4_out7_real(Stage4_out7_real),
	.Stage4_out7_imag(Stage4_out7_imag),
	.Stage4_out8_real(Stage4_out8_real),
	.Stage4_out8_imag(Stage4_out8_imag),
	.Stage4_out9_real(Stage4_out9_real),
	.Stage4_out9_imag(Stage4_out9_imag),
	.Stage4_out10_real(Stage4_out10_real),
	.Stage4_out10_imag(Stage4_out10_imag),
	.Stage4_out11_real(Stage4_out11_real),
	.Stage4_out11_imag(Stage4_out11_imag),
	.Stage4_out12_real(Stage4_out12_real),
	.Stage4_out12_imag(Stage4_out12_imag),
	.Stage4_out13_real(Stage4_out13_real),
	.Stage4_out13_imag(Stage4_out13_imag),
	.Stage4_out14_real(Stage4_out14_real),
	.Stage4_out14_imag(Stage4_out14_imag),
	.Stage4_out15_real(Stage4_out15_real),
	.Stage4_out15_imag(Stage4_out15_imag),
	.Stage4_out16_real(Stage4_out16_real),
	.Stage4_out16_imag(Stage4_out16_imag),
	.Stage4_out17_real(Stage4_out17_real),
	.Stage4_out17_imag(Stage4_out17_imag),
	.Stage4_out18_real(Stage4_out18_real),
	.Stage4_out18_imag(Stage4_out18_imag),
	.Stage4_out19_real(Stage4_out19_real),
	.Stage4_out19_imag(Stage4_out19_imag),
	.Stage4_out20_real(Stage4_out20_real),
	.Stage4_out20_imag(Stage4_out20_imag),
	.Stage4_out21_real(Stage4_out21_real),
	.Stage4_out21_imag(Stage4_out21_imag),
	.Stage4_out22_real(Stage4_out22_real),
	.Stage4_out22_imag(Stage4_out22_imag),
	.Stage4_out23_real(Stage4_out23_real),
	.Stage4_out23_imag(Stage4_out23_imag),
	.Stage4_out24_real(Stage4_out24_real),
	.Stage4_out24_imag(Stage4_out24_imag),
	.Stage4_out25_real(Stage4_out25_real),
	.Stage4_out25_imag(Stage4_out25_imag),
	.Stage4_out26_real(Stage4_out26_real),
	.Stage4_out26_imag(Stage4_out26_imag),
	.Stage4_out27_real(Stage4_out27_real),
	.Stage4_out27_imag(Stage4_out27_imag),
	.Stage4_out28_real(Stage4_out28_real),
	.Stage4_out28_imag(Stage4_out28_imag),
	.Stage4_out29_real(Stage4_out29_real),
	.Stage4_out29_imag(Stage4_out29_imag),
	.Stage4_out30_real(Stage4_out30_real),
	.Stage4_out30_imag(Stage4_out30_imag),
	.Stage4_out31_real(Stage4_out31_real),
	.Stage4_out31_imag(Stage4_out31_imag),
	.Stage5_out0_real(FFT_RESULT_0_real),
	.Stage5_out0_imag(FFT_RESULT_0_imag),
	.Stage5_out1_real(FFT_RESULT_1_real),
	.Stage5_out1_imag(FFT_RESULT_1_imag),
	.Stage5_out2_real(FFT_RESULT_2_real),
	.Stage5_out2_imag(FFT_RESULT_2_imag),
	.Stage5_out3_real(FFT_RESULT_3_real),
	.Stage5_out3_imag(FFT_RESULT_3_imag),
	.Stage5_out4_real(FFT_RESULT_4_real),
	.Stage5_out4_imag(FFT_RESULT_4_imag),
	.Stage5_out5_real(FFT_RESULT_5_real),
	.Stage5_out5_imag(FFT_RESULT_5_imag),
	.Stage5_out6_real(FFT_RESULT_6_real),
	.Stage5_out6_imag(FFT_RESULT_6_imag),
	.Stage5_out7_real(FFT_RESULT_7_real),
	.Stage5_out7_imag(FFT_RESULT_7_imag),
	.Stage5_out8_real(FFT_RESULT_8_real),
	.Stage5_out8_imag(FFT_RESULT_8_imag),
	.Stage5_out9_real(FFT_RESULT_9_real),
	.Stage5_out9_imag(FFT_RESULT_9_imag),
	.Stage5_out10_real(FFT_RESULT_10_real),
	.Stage5_out10_imag(FFT_RESULT_10_imag),
	.Stage5_out11_real(FFT_RESULT_11_real),
	.Stage5_out11_imag(FFT_RESULT_11_imag),
	.Stage5_out12_real(FFT_RESULT_12_real),
	.Stage5_out12_imag(FFT_RESULT_12_imag),
	.Stage5_out13_real(FFT_RESULT_13_real),
	.Stage5_out13_imag(FFT_RESULT_13_imag),
	.Stage5_out14_real(FFT_RESULT_14_real),
	.Stage5_out14_imag(FFT_RESULT_14_imag),
	.Stage5_out15_real(FFT_RESULT_15_real),
	.Stage5_out15_imag(FFT_RESULT_15_imag),
	.Stage5_out16_real(FFT_RESULT_16_real),
	.Stage5_out16_imag(FFT_RESULT_16_imag),
	.Stage5_out17_real(FFT_RESULT_17_real),
	.Stage5_out17_imag(FFT_RESULT_17_imag),
	.Stage5_out18_real(FFT_RESULT_18_real),
	.Stage5_out18_imag(FFT_RESULT_18_imag),
	.Stage5_out19_real(FFT_RESULT_19_real),
	.Stage5_out19_imag(FFT_RESULT_19_imag),
	.Stage5_out20_real(FFT_RESULT_20_real),
	.Stage5_out20_imag(FFT_RESULT_20_imag),
	.Stage5_out21_real(FFT_RESULT_21_real),
	.Stage5_out21_imag(FFT_RESULT_21_imag),
	.Stage5_out22_real(FFT_RESULT_22_real),
	.Stage5_out22_imag(FFT_RESULT_22_imag),
	.Stage5_out23_real(FFT_RESULT_23_real),
	.Stage5_out23_imag(FFT_RESULT_23_imag),
	.Stage5_out24_real(FFT_RESULT_24_real),
	.Stage5_out24_imag(FFT_RESULT_24_imag),
	.Stage5_out25_real(FFT_RESULT_25_real),
	.Stage5_out25_imag(FFT_RESULT_25_imag),
	.Stage5_out26_real(FFT_RESULT_26_real),
	.Stage5_out26_imag(FFT_RESULT_26_imag),
	.Stage5_out27_real(FFT_RESULT_27_real),
	.Stage5_out27_imag(FFT_RESULT_27_imag),
	.Stage5_out28_real(FFT_RESULT_28_real),
	.Stage5_out28_imag(FFT_RESULT_28_imag),
	.Stage5_out29_real(FFT_RESULT_29_real),
	.Stage5_out29_imag(FFT_RESULT_29_imag),
	.Stage5_out30_real(FFT_RESULT_30_real),
	.Stage5_out30_imag(FFT_RESULT_30_imag),
	.Stage5_out31_real(FFT_RESULT_31_real),
	.Stage5_out31_imag(FFT_RESULT_31_imag),
	.Constant_W0_real(Constant_W0_real),
	.Constant_W0_imag(Constant_W0_imag),
	.Constant_W1_real(Constant_W1_real),
	.Constant_W1_imag(Constant_W1_imag),
	.Constant_W2_real(Constant_W2_real),
	.Constant_W2_imag(Constant_W2_imag),
	.Constant_W3_real(Constant_W3_real),
	.Constant_W3_imag(Constant_W3_imag),
	.Constant_W4_real(Constant_W4_real),
	.Constant_W4_imag(Constant_W4_imag),
	.Constant_W5_real(Constant_W5_real),
	.Constant_W5_imag(Constant_W5_imag),
	.Constant_W6_real(Constant_W6_real),
	.Constant_W6_imag(Constant_W6_imag),
	.Constant_W7_real(Constant_W7_real),
	.Constant_W7_imag(Constant_W7_imag),
	.Constant_W8_real(Constant_W8_real),
	.Constant_W8_imag(Constant_W8_imag),
	.Constant_W9_real(Constant_W9_real),
	.Constant_W9_imag(Constant_W9_imag),
	.Constant_W10_real(Constant_W10_real),
	.Constant_W10_imag(Constant_W10_imag),
	.Constant_W11_real(Constant_W11_real),
	.Constant_W11_imag(Constant_W11_imag),
	.Constant_W12_real(Constant_W12_real),
	.Constant_W12_imag(Constant_W12_imag),
	.Constant_W13_real(Constant_W13_real),
	.Constant_W13_imag(Constant_W13_imag),
	.Constant_W14_real(Constant_W14_real),
	.Constant_W14_imag(Constant_W14_imag),
	.Constant_W15_real(Constant_W15_real),
	.Constant_W15_imag(Constant_W15_imag)
);



endmodule